`ifndef PARAMETER_H_
`define PARAMETER_H_

// Parameter file for RISC processor
`define col 16
`define row_i 15
`define row_d 8
`define filename "./test/50001111_50001212.o"
`define simulation_time #160

`endif
